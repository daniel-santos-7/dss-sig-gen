
library IEEE;
use IEEE.std_logic_1164.all;

package sine_lut_pkg is
    
    constant LUT_ADDR_BITS : natural := 8;

    constant OUT_RES_BITS  : natural := 12;

    type sine_lut_array is array (0 to 2 ** LUT_ADDR_BITS-1) of std_logic_vector(OUT_RES_BITS-1 downto 0);

    constant SINE_TABLE : sine_lut_array := (
        x"000",
		x"000",
		x"000",
		x"001",
		x"002",
		x"003",
		x"005",
		x"007",
		x"009",
		x"00c",
		x"00f",
		x"012",
		x"016",
		x"019",
		x"01e",
		x"022",
		x"027",
		x"02c",
		x"031",
		x"037",
		x"03d",
		x"043",
		x"04a",
		x"050",
		x"058",
		x"05f",
		x"067",
		x"06f",
		x"077",
		x"080",
		x"089",
		x"092",
		x"09b",
		x"0a5",
		x"0af",
		x"0b9",
		x"0c4",
		x"0cf",
		x"0da",
		x"0e6",
		x"0f1",
		x"0fd",
		x"109",
		x"116",
		x"123",
		x"130",
		x"13d",
		x"14b",
		x"158",
		x"167",
		x"175",
		x"183",
		x"192",
		x"1a1",
		x"1b1",
		x"1c0",
		x"1d0",
		x"1e0",
		x"1f0",
		x"201",
		x"212",
		x"223",
		x"234",
		x"245",
		x"257",
		x"269",
		x"27b",
		x"28d",
		x"2a0",
		x"2b3",
		x"2c5",
		x"2d9",
		x"2ec",
		x"2ff",
		x"313",
		x"327",
		x"33b",
		x"34f",
		x"364",
		x"378",
		x"38d",
		x"3a2",
		x"3b7",
		x"3cd",
		x"3e2",
		x"3f8",
		x"40e",
		x"423",
		x"43a",
		x"450",
		x"466",
		x"47d",
		x"493",
		x"4aa",
		x"4c1",
		x"4d8",
		x"4ef",
		x"506",
		x"51e",
		x"535",
		x"54d",
		x"565",
		x"57c",
		x"594",
		x"5ac",
		x"5c4",
		x"5dd",
		x"5f5",
		x"60d",
		x"626",
		x"63e",
		x"657",
		x"66f",
		x"688",
		x"6a1",
		x"6b9",
		x"6d2",
		x"6eb",
		x"704",
		x"71d",
		x"736",
		x"74f",
		x"768",
		x"781",
		x"79a",
		x"7b3",
		x"7cc",
		x"7e5",
		x"7ff",
		x"818",
		x"831",
		x"84a",
		x"863",
		x"87c",
		x"895",
		x"8ae",
		x"8c7",
		x"8e0",
		x"8f9",
		x"912",
		x"92b",
		x"944",
		x"95c",
		x"975",
		x"98e",
		x"9a6",
		x"9bf",
		x"9d7",
		x"9f0",
		x"a08",
		x"a20",
		x"a39",
		x"a51",
		x"a69",
		x"a81",
		x"a98",
		x"ab0",
		x"ac8",
		x"adf",
		x"af7",
		x"b0e",
		x"b25",
		x"b3c",
		x"b53",
		x"b6a",
		x"b80",
		x"b97",
		x"bad",
		x"bc3",
		x"bda",
		x"bef",
		x"c05",
		x"c1b",
		x"c30",
		x"c46",
		x"c5b",
		x"c70",
		x"c85",
		x"c99",
		x"cae",
		x"cc2",
		x"cd6",
		x"cea",
		x"cfe",
		x"d11",
		x"d24",
		x"d38",
		x"d4a",
		x"d5d",
		x"d70",
		x"d82",
		x"d94",
		x"da6",
		x"db8",
		x"dc9",
		x"dda",
		x"deb",
		x"dfc",
		x"e0d",
		x"e1d",
		x"e2d",
		x"e3d",
		x"e4c",
		x"e5c",
		x"e6b",
		x"e7a",
		x"e88",
		x"e96",
		x"ea5",
		x"eb2",
		x"ec0",
		x"ecd",
		x"eda",
		x"ee7",
		x"ef4",
		x"f00",
		x"f0c",
		x"f17",
		x"f23",
		x"f2e",
		x"f39",
		x"f44",
		x"f4e",
		x"f58",
		x"f62",
		x"f6b",
		x"f74",
		x"f7d",
		x"f86",
		x"f8e",
		x"f96",
		x"f9e",
		x"fa5",
		x"fad",
		x"fb3",
		x"fba",
		x"fc0",
		x"fc6",
		x"fcc",
		x"fd1",
		x"fd6",
		x"fdb",
		x"fdf",
		x"fe4",
		x"fe7",
		x"feb",
		x"fee",
		x"ff1",
		x"ff4",
		x"ff6",
		x"ff8",
		x"ffa",
		x"ffb",
		x"ffc",
		x"ffd",
		x"ffd"
    );

end package sine_lut_pkg;
    
