library IEEE;
use IEEE.std_logic_1164.all;

package sine_lut_pkg is
    
    constant LUT_ADDR_BITS : natural := 8;

    constant OUT_RES_BITS  : natural := 12;

    type sine_lut_array is array (0 to 2 ** LUT_ADDR_BITS-1) of std_logic_vector(OUT_RES_BITS-1 downto 0);

    constant SINE_TABLE : sine_lut_array := (
        x"801",
		x"802",
		x"802",
		x"803",
		x"804",
		x"805",
		x"807",
		x"809",
		x"80b",
		x"80e",
		x"811",
		x"814",
		x"818",
		x"81b",
		x"820",
		x"824",
		x"829",
		x"82e",
		x"833",
		x"839",
		x"83f",
		x"845",
		x"84c",
		x"852",
		x"85a",
		x"861",
		x"869",
		x"871",
		x"879",
		x"882",
		x"88b",
		x"894",
		x"89d",
		x"8a7",
		x"8b1",
		x"8bb",
		x"8c6",
		x"8d1",
		x"8dc",
		x"8e8",
		x"8f3",
		x"8ff",
		x"90b",
		x"918",
		x"925",
		x"932",
		x"93f",
		x"94d",
		x"95a",
		x"969",
		x"977",
		x"985",
		x"994",
		x"9a3",
		x"9b3",
		x"9c2",
		x"9d2",
		x"9e2",
		x"9f2",
		x"a03",
		x"a14",
		x"a25",
		x"a36",
		x"a47",
		x"a59",
		x"a6b",
		x"a7d",
		x"a8f",
		x"aa2",
		x"ab5",
		x"ac7",
		x"adb",
		x"aee",
		x"b01",
		x"b15",
		x"b29",
		x"b3d",
		x"b51",
		x"b66",
		x"b7a",
		x"b8f",
		x"ba4",
		x"bb9",
		x"bcf",
		x"be4",
		x"bfa",
		x"c10",
		x"c25",
		x"c3c",
		x"c52",
		x"c68",
		x"c7f",
		x"c95",
		x"cac",
		x"cc3",
		x"cda",
		x"cf1",
		x"d08",
		x"d20",
		x"d37",
		x"d4f",
		x"d67",
		x"d7e",
		x"d96",
		x"dae",
		x"dc6",
		x"ddf",
		x"df7",
		x"e0f",
		x"e28",
		x"e40",
		x"e59",
		x"e71",
		x"e8a",
		x"ea3",
		x"ebb",
		x"ed4",
		x"eed",
		x"f06",
		x"f1f",
		x"f38",
		x"f51",
		x"f6a",
		x"f83",
		x"f9c",
		x"fb5",
		x"fce",
		x"fe7",
		x"000",
		x"019",
		x"032",
		x"04b",
		x"064",
		x"07d",
		x"096",
		x"0af",
		x"0c8",
		x"0e1",
		x"0fa",
		x"113",
		x"12c",
		x"145",
		x"15d",
		x"176",
		x"18f",
		x"1a7",
		x"1c0",
		x"1d8",
		x"1f1",
		x"209",
		x"221",
		x"23a",
		x"252",
		x"26a",
		x"282",
		x"299",
		x"2b1",
		x"2c9",
		x"2e0",
		x"2f8",
		x"30f",
		x"326",
		x"33d",
		x"354",
		x"36b",
		x"381",
		x"398",
		x"3ae",
		x"3c4",
		x"3db",
		x"3f0",
		x"406",
		x"41c",
		x"431",
		x"447",
		x"45c",
		x"471",
		x"486",
		x"49a",
		x"4af",
		x"4c3",
		x"4d7",
		x"4eb",
		x"4ff",
		x"512",
		x"525",
		x"539",
		x"54b",
		x"55e",
		x"571",
		x"583",
		x"595",
		x"5a7",
		x"5b9",
		x"5ca",
		x"5db",
		x"5ec",
		x"5fd",
		x"60e",
		x"61e",
		x"62e",
		x"63e",
		x"64d",
		x"65d",
		x"66c",
		x"67b",
		x"689",
		x"697",
		x"6a6",
		x"6b3",
		x"6c1",
		x"6ce",
		x"6db",
		x"6e8",
		x"6f5",
		x"701",
		x"70d",
		x"718",
		x"724",
		x"72f",
		x"73a",
		x"745",
		x"74f",
		x"759",
		x"763",
		x"76c",
		x"775",
		x"77e",
		x"787",
		x"78f",
		x"797",
		x"79f",
		x"7a6",
		x"7ae",
		x"7b4",
		x"7bb",
		x"7c1",
		x"7c7",
		x"7cd",
		x"7d2",
		x"7d7",
		x"7dc",
		x"7e0",
		x"7e5",
		x"7e8",
		x"7ec",
		x"7ef",
		x"7f2",
		x"7f5",
		x"7f7",
		x"7f9",
		x"7fb",
		x"7fc",
		x"7fd",
		x"7fe",
		x"7fe"
    );

end package sine_lut_pkg;
