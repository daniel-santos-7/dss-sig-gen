library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity sine_lut is
    generic (
        LUT_ADDR_BITS : natural := 8;
        OUT_RES_BITS  : natural := 12
    );
    port (
        rst_n : in  std_logic;
        clk   : in  std_logic;
        addr  : in  std_logic_vector(LUT_ADDR_BITS-1 downto 0);
        wave  : out std_logic_vector(OUT_RES_BITS-1 downto 0)
    );
end entity sine_lut;

architecture rtl of sine_lut is

    type sine_lut_array is array (natural range 0 to 255) of std_logic_vector(11 downto 0);

    constant SINE_TABLE : sine_lut_array := (
        X"000",
        X"019",
        X"032",
        X"04B",
        X"064",
        X"07D",
        X"096",
        X"0AF",
        X"0C8",
        X"0E2",
        X"0FB",
        X"114",
        X"12D",
        X"146",
        X"15F",
        X"178",
        X"191",
        X"1AA",
        X"1C3",
        X"1DC",
        X"1F5",
        X"20E",
        X"227",
        X"23F",
        X"258",
        X"271",
        X"28A",
        X"2A3",
        X"2BC",
        X"2D4",
        X"2ED",
        X"306",
        X"31E",
        X"337",
        X"350",
        X"368",
        X"381",
        X"399",
        X"3B2",
        X"3CA",
        X"3E3",
        X"3FB",
        X"413",
        X"42B",
        X"444",
        X"45C",
        X"474",
        X"48C",
        X"4A4",
        X"4BC",
        X"4D4",
        X"4EC",
        X"504",
        X"51C",
        X"534",
        X"54B",
        X"563",
        X"57B",
        X"592",
        X"5AA",
        X"5C1",
        X"5D9",
        X"5F0",
        X"607",
        X"61F",
        X"636",
        X"64D",
        X"664",
        X"67B",
        X"692",
        X"6A9",
        X"6C0",
        X"6D6",
        X"6ED",
        X"704",
        X"71A",
        X"731",
        X"747",
        X"75D",
        X"774",
        X"78A",
        X"7A0",
        X"7B6",
        X"7CC",
        X"7E2",
        X"7F8",
        X"80D",
        X"823",
        X"839",
        X"84E",
        X"864",
        X"879",
        X"88E",
        X"8A4",
        X"8B9",
        X"8CE",
        X"8E3",
        X"8F7",
        X"90C",
        X"921",
        X"935",
        X"94A",
        X"95E",
        X"973",
        X"987",
        X"99B",
        X"9AF",
        X"9C3",
        X"9D7",
        X"9EB",
        X"9FE",
        X"A12",
        X"A25",
        X"A39",
        X"A4C",
        X"A5F",
        X"A72",
        X"A85",
        X"A98",
        X"AAB",
        X"ABE",
        X"AD0",
        X"AE3",
        X"AF5",
        X"B07",
        X"B19",
        X"B2B",
        X"B3D",
        X"B4F",
        X"B61",
        X"B72",
        X"B84",
        X"B95",
        X"BA7",
        X"BB8",
        X"BC9",
        X"BDA",
        X"BEB",
        X"BFB",
        X"C0C",
        X"C1C",
        X"C2D",
        X"C3D",
        X"C4D",
        X"C5D",
        X"C6D",
        X"C7D",
        X"C8C",
        X"C9C",
        X"CAB",
        X"CBA",
        X"CCA",
        X"CD9",
        X"CE8",
        X"CF6",
        X"D05",
        X"D14",
        X"D22",
        X"D30",
        X"D3E",
        X"D4C",
        X"D5A",
        X"D68",
        X"D76",
        X"D83",
        X"D91",
        X"D9E",
        X"DAB",
        X"DB8",
        X"DC5",
        X"DD1",
        X"DDE",
        X"DEB",
        X"DF7",
        X"E03",
        X"E0F",
        X"E1B",
        X"E27",
        X"E32",
        X"E3E",
        X"E49",
        X"E54",
        X"E60",
        X"E6B",
        X"E75",
        X"E80",
        X"E8B",
        X"E95",
        X"E9F",
        X"EA9",
        X"EB3",
        X"EBD",
        X"EC7",
        X"ED0",
        X"EDA",
        X"EE3",
        X"EEC",
        X"EF5",
        X"EFE",
        X"F07",
        X"F0F",
        X"F18",
        X"F20",
        X"F28",
        X"F30",
        X"F38",
        X"F3F",
        X"F47",
        X"F4E",
        X"F55",
        X"F5C",
        X"F63",
        X"F6A",
        X"F71",
        X"F77",
        X"F7E",
        X"F84",
        X"F8A",
        X"F90",
        X"F95",
        X"F9B",
        X"FA0",
        X"FA6",
        X"FAB",
        X"FB0",
        X"FB5",
        X"FB9",
        X"FBE",
        X"FC2",
        X"FC6",
        X"FCA",
        X"FCE",
        X"FD2",
        X"FD6",
        X"FD9",
        X"FDD",
        X"FE0",
        X"FE3",
        X"FE6",
        X"FE8",
        X"FEB",
        X"FED",
        X"FEF",
        X"FF1",
        X"FF3",
        X"FF5",
        X"FF7",
        X"FF8",
        X"FFA",
        X"FFB",
        X"FFC",
        X"FFD",
        X"FFD",
        X"FFE",
        X"FFE",
        X"FFE"
    );

    signal wave_reg : std_logic_vector(OUT_RES_BITS-1 downto 0);

begin

    wave_reg_logic : process(rst_n, clk)
        variable idx : natural range 0 to 255;
    begin
        if rising_edge(clk) then
            if rst_n = '0' then
                wave_reg <= (others => '0');
            else
                idx := to_integer(unsigned(addr));
                wave_reg <= SINE_TABLE(idx);
            end if ;
        end if ;
    end process ; -- wave_reg_logic

    -- Assign register to output
    wave <= wave_reg;

end architecture rtl;