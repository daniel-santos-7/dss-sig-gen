library IEEE;
use IEEE.std_logic_1164.all;

package sine_lut_pkg is
    
    constant LUT_ADDR_BITS : natural := 8;

    constant OUT_RES_BITS  : natural := 12;

    type sine_lut_array is array (0 to 2 ** LUT_ADDR_BITS-1) of std_logic_vector(OUT_RES_BITS-1 downto 0);

    constant SINE_TABLE : sine_lut_array := (
		x"000",
		x"00c",
		x"019",
		x"025",
		x"032",
		x"03e",
		x"04b",
		x"057",
		x"064",
		x"070",
		x"07d",
		x"08a",
		x"096",
		x"0a3",
		x"0af",
		x"0bc",
		x"0c8",
		x"0d5",
		x"0e1",
		x"0ee",
		x"0fa",
		x"107",
		x"113",
		x"11f",
		x"12c",
		x"138",
		x"145",
		x"151",
		x"15d",
		x"16a",
		x"176",
		x"183",
		x"18f",
		x"19b",
		x"1a7",
		x"1b4",
		x"1c0",
		x"1cc",
		x"1d8",
		x"1e5",
		x"1f1",
		x"1fd",
		x"209",
		x"215",
		x"221",
		x"22e",
		x"23a",
		x"246",
		x"252",
		x"25e",
		x"26a",
		x"276",
		x"282",
		x"28e",
		x"299",
		x"2a5",
		x"2b1",
		x"2bd",
		x"2c9",
		x"2d4",
		x"2e0",
		x"2ec",
		x"2f8",
		x"303",
		x"30f",
		x"31a",
		x"326",
		x"332",
		x"33d",
		x"348",
		x"354",
		x"35f",
		x"36b",
		x"376",
		x"381",
		x"38d",
		x"398",
		x"3a3",
		x"3ae",
		x"3b9",
		x"3c4",
		x"3d0",
		x"3db",
		x"3e6",
		x"3f0",
		x"3fb",
		x"406",
		x"411",
		x"41c",
		x"427",
		x"431",
		x"43c",
		x"447",
		x"451",
		x"45c",
		x"466",
		x"471",
		x"47b",
		x"486",
		x"490",
		x"49a",
		x"4a4",
		x"4af",
		x"4b9",
		x"4c3",
		x"4cd",
		x"4d7",
		x"4e1",
		x"4eb",
		x"4f5",
		x"4ff",
		x"508",
		x"512",
		x"51c",
		x"525",
		x"52f",
		x"539",
		x"542",
		x"54b",
		x"555",
		x"55e",
		x"567",
		x"571",
		x"57a",
		x"583",
		x"58c",
		x"595",
		x"59e",
		x"5a7",
		x"5b0",
		x"5b9",
		x"5c1",
		x"5ca",
		x"5d3",
		x"5db",
		x"5e4",
		x"5ec",
		x"5f5",
		x"5fd",
		x"605",
		x"60e",
		x"616",
		x"61e",
		x"626",
		x"62e",
		x"636",
		x"63e",
		x"645",
		x"64d",
		x"655",
		x"65d",
		x"664",
		x"66c",
		x"673",
		x"67b",
		x"682",
		x"689",
		x"690",
		x"697",
		x"69f",
		x"6a6",
		x"6ac",
		x"6b3",
		x"6ba",
		x"6c1",
		x"6c8",
		x"6ce",
		x"6d5",
		x"6db",
		x"6e2",
		x"6e8",
		x"6ee",
		x"6f5",
		x"6fb",
		x"701",
		x"707",
		x"70d",
		x"713",
		x"718",
		x"71e",
		x"724",
		x"72a",
		x"72f",
		x"735",
		x"73a",
		x"73f",
		x"745",
		x"74a",
		x"74f",
		x"754",
		x"759",
		x"75e",
		x"763",
		x"767",
		x"76c",
		x"771",
		x"775",
		x"77a",
		x"77e",
		x"783",
		x"787",
		x"78b",
		x"78f",
		x"793",
		x"797",
		x"79b",
		x"79f",
		x"7a3",
		x"7a6",
		x"7aa",
		x"7ae",
		x"7b1",
		x"7b4",
		x"7b8",
		x"7bb",
		x"7be",
		x"7c1",
		x"7c4",
		x"7c7",
		x"7ca",
		x"7cd",
		x"7cf",
		x"7d2",
		x"7d5",
		x"7d7",
		x"7da",
		x"7dc",
		x"7de",
		x"7e0",
		x"7e2",
		x"7e5",
		x"7e6",
		x"7e8",
		x"7ea",
		x"7ec",
		x"7ee",
		x"7ef",
		x"7f1",
		x"7f2",
		x"7f3",
		x"7f5",
		x"7f6",
		x"7f7",
		x"7f8",
		x"7f9",
		x"7fa",
		x"7fb",
		x"7fb",
		x"7fc",
		x"7fd",
		x"7fd",
		x"7fe",
		x"7fe",
		x"7fe",
		x"7fe",
		x"7fe"
	);

end package sine_lut_pkg;
